typedef struct packed {
    logic [7:0] port0_count;
    logic [7:0] port1_count;
    logic [7:0] port2_count;
} config_t;

